module memory (
    input i_Clk,
    input i_Rst,
    input [7:0] i_Data,
    input i_Loa
);
    
endmodule
module sleep(
    input i_Clk,            // Input Clock
    input i_Start,          // Start Sleep
    output o_Done          // Output data bus
);
    reg 

endmodule